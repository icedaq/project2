localparam [31:0] biases [9 : 0] = {32'h000000c3, 32'h00000149, 32'h0000011c, 32'h000000d9, 32'h0000010b, 32'h000001fa, 32'h000000f9, 32'h0000017c, 32'h00000000, 32'h000000de}